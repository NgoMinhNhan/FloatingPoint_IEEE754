`include "chia.v"
module chia_tb;
	reg [31:0]A,B;
	wire [31:0]KQ;
	chia abcd(.a(A[31:0]),.b(B[31:0]),.result(KQ[31:0]));
	initial begin
/*---------------------------------------------------------------*/
	#0	B=32'b0_01111111_10000000000000000000000;
	A=32'b0_01111111_10000000000000000000000;
	#10     A=32'b01111111111111111111111111111111; //NaN
		B=32'b01111111111111111111111111111111; //NaN	
	#10	B=32'b00000000000000000000000000000000; //+Zero
	#10	B=32'b10000000000000000000000000000000; //-Zero
	#10	B=32'b01111111100000000000000000000000; //+Inf
	#10	B=32'b11111111100000000000000000000000; //-Inf
	#10	B=32'b01000001010001011000011110010100;//+12.3456
	#10	B=32'b11000001010001011000011110010100;//-12.3456
	#10

	
	B=32'b1_01111110_00000000000000000000000;
	A=32'b1_10000000_01000000000000000000000;
	#100
	B=32'b0_01111110_00000000000000000000000;
	A=32'b0_01111110_00000000000000000000000;
	#100;
	end
	
initial begin

$vcdplusfile ("chia.vpd");
$vcdpluson ();
end
endmodule
`include "power.v"
module power_tb();

reg [31:0] base;
reg [31:0] exp;

wire [31:0] out;


power power_A_B(.a_base(base),.b_exp(exp), .result(out));

initial begin
	
	#10
	base = 32'b01000100011110100000000000000000; // 1000
	exp  = 32'b01000000101000000000000000000000; // 5
	 #10
	 base = 32'b01000000110000000000000000000000; // 6
	 exp  = 32'b01000001000100000000000000000000; // 9
	 #10
	 base = 32'b00111110110000000000000000000000; // 0.375
	 exp  = 32'b00111110110011001100110011001101; // 0.4
	 #10
	 base = 32'b00111110110011001100110011001101; // 0.4
	 exp  = 32'b00111110110011001100110011001101; // 0.4
	 #10
	 base = 32'b00111110010011001100110011001101; // 0.2
	 exp  = 32'b00111110110011001100110011001101; // 0.4
	
end

endmodule 
initial begin
$vcdplusfile ("nth_root_tb.vpd");
$vcdpluson ();
end
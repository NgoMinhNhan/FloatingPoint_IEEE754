module nhan_tb;
	reg [31:0]A,B;
	wire [31:0]result;	
	
	nhan m7(.a(A[31:0]),.b(B[31:0]),.result(result[31:0]));
	initial begin
	#0	

	A=32'b0_01111111_00000000000000000000000; //1
	B=32'b0_01111111_00000000000000000000000; //1
        #10
A=32'b1100_1011_1111_1111_1001_0101_1011_0000; 
B=32'b1101_0000_0000_1111_0000_1101_0001_1000;
       
       #10	

	A=32'b0_01111111_00000000000000000000000; //0.02345
	B=32'b0_01111010_00011011000111011001001; //0.03456
#10	
	A=32'b0_01111111_10000000000000000000000; //0.02345
	B=32'b0_01111111_11000000000000000000000; //0.03456

#10
	A=32'b0_11111111_11000000000000000000000;
	B=32'b0_11111111_10000000000000000000000;
	#10
	A=32'b0_00000001_11000000000000000000000;
	B=32'b1_00000001_00000000000000000000000;
	#10
	A=32'b0_11111110_11000000000000000000000;	// ex(A) + ex(B) -127 = 8'b 1111_1111
	B=32'b1_10000000_00000000000000000000000;
	#10
	A=32'b1_11111110_11111111111111111111111;
	B=32'b0_00000001_11111111111111111111111;
	#10
	A=32'b1_00000000_11000000000000000000011;
	B=32'b1_00000000_11000000000000000000011;
	#10
	A=32'b1_00000001_11000000000000000000000;
	B=32'b1_00000010_11000000000000000000000;
	#10
	A=32'b0_10000000_00101100001010001111011; // 2.345
	B=32'b0_10000000_10111010010111100011011; // 3.456
	
	#100
	;
end

initial begin
$vcdplusflie ("nhan_tb.vpd")
$vcdpluson ();
end
endmodule